`timescale 1ns / 1ns

module D-Flop(
    );


endmodule
